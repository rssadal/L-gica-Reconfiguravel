LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;


ENTITY PROJETO IS
	PORT(
		
		ENTRADA_1: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		SINAL_1: IN STD_LOGIC;
		ENTRADA_2: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		SINAL_2: IN STD_LOGIC;		

		RESULTADO_DISPLAY_1: OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
		RESULTADO_DISPLAY_2: OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
		RESULTADO_DISPLAY_3: OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
		RESULTADO_LEDS: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		
		SAIDA_OPERACAO_DISPLAY: OUT STD_LOGIC_VECTOR (0 TO 6);	
		
		PUSH_RESULTADO: IN STD_LOGIC;
		PUSH_OPERACAO: IN STD_LOGIC;
		RESET: IN STD_LOGIC;
		CLOCK: IN STD_LOGIC;
		LED_REFERENCIA: OUT STD_LOGIC
		
	);
END PROJETO;

ARCHITECTURE MODELO OF PROJETO IS 

CONSTANT CLOCK_FREE : INTEGER := 50e6;
SIGNAL TICKS : INTEGER := 0;
SIGNAL SEGUNDOS: INTEGER := 0;

SIGNAL OPERACAO: INTEGER := 1;

-- GUARDANDO RESULTADOS
SIGNAL RESULTADO_ARI: INTEGER := 0;
SIGNAL RESULTADO_LOG: STD_LOGIC_VECTOR (3 DOWNTO 0);

-- TRANSFORMANDO ENTRADA EM VALOR NÚMERICO
SIGNAL VALOR_1: INTEGER := TO_INTEGER(UNSIGNED(ENTRADA_1)); 
SIGNAL VALOR_2: INTEGER := TO_INTEGER(UNSIGNED(ENTRADA_2));


BEGIN
	
	PROCESS (CLOCK) IS
	BEGIN
	
		IF RISING_EDGE(CLOCK) THEN -- NA BORDA DO CLOCK
			IF TICKS = CLOCK_FREE - 1 THEN
				TICKS <= 0;
				-- CONTADOR DE TICKS
				IF SEGUNDOS = 3 THEN -- VAI aGIR APENAS QUANDO BATER 3S 
					SEGUNDOS <= 0;
					LED_REFERENCIA <= '1';
					CASE OPERACAO IS
						
						WHEN 1 => -- SOMA
						
							IF SINAL_1 = '0' THEN
								 VALOR_1 <= -VALOR_1;
							END IF;
							IF SINAL_2 = '0' THEN
								 VALOR_2 <= -VALOR_2;
							END IF;
							
							RESULTADO_ARI <= VALOR_1 + VALOR_2;
							
						WHEN 2 => -- ADIÇÃO
							
							IF SINAL_1 = '0' THEN
								 VALOR_1 <= -VALOR_1;
							END IF;
							IF SINAL_2 = '0' THEN
								 VALOR_2 <= -VALOR_2;
							END IF;
							
							RESULTADO_ARI <= VALOR_1 - VALOR_2;
						
						WHEN 3 => -- E
							
							RESULTADO_LOG <= ENTRADA_1 AND ENTRADA_2;
							
						WHEN 4 => -- OU
							
							RESULTADO_LOG <= ENTRADA_1 OR ENTRADA_2;
							
						WHEN 5 => -- OU EXCLUSUVIO
							
							RESULTADO_LOG <= ENTRADA_1 XOR ENTRADA_2;
							
						WHEN OTHERS => -- COMPLEMENTO	
							 
							RESULTADO_LOG <= NOT ENTRADA_1;
							
					END CASE;
					
				ELSE
					SEGUNDOS <= SEGUNDOS + 1;
					LED_REFERENCIA <= '0';
				END IF;
				
			ELSE
				TICKS <= ticks + 1;
			END IF;
		END IF;
		
		IF RESET = '0' THEN -- RESETA TUDO E APAGA O DISPLAY
			TICKS <= 0;
			SEGUNDOS <= 0;
			OPERACAO <= 1;
			SAIDA_RESULTADO <= "1111111";
			LED_REFERENCIA <= '1';
			-- RESETAR TUDO 
		END IF;
		
		IF PUSH_OPERACAO = '0' THEN -- INCREMENTO DA OPERAÇÃO
			OPERACAO <= OPERACAO + 1;
			IF OPERACAO = 6 THEN
				OPERACAO <= 1;
			END IF;
		END IF;
		
		IF PUSH_RESULTADO = '0' THEN -- MOSTRAR O RESULTADO
			IF OPERACAO < 3 THEN
					-- OPERAÇÕES ARITMETICAS
			ELSE
			      -- OPERAÇÕES LÓGICAS
			END IF;
		END IF;
										 
		SAIDA_OPERACAO_DISPLAY <=
        "1001111" WHEN OPERACAO = 1, -- '1'
        "0010010" WHEN OPERACAO = 2, -- '2'
        "0000110" WHEN OPERACAO = 3, -- '3'
        "1001100" WHEN OPERACAO = 4, -- '4'
        "0100100" WHEN OPERACAO = 5, -- '5'
        "0100000" WHEN OTHERS;       -- '6'
		
	END PROCESS;

END MODELO;