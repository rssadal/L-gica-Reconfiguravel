LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;


ENTITY PROJETO IS
	PORT(
		
		ENTRADA_1: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		SINAL_1: IN STD_LOGIC;
		ENTRADA_2: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		SINAL_2: IN STD_LOGIC;		

		RESULTADO_DISPLAY_1: OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
		RESULTADO_DISPLAY_2: OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
		RESULTADO_DISPLAY_3: OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
		RESULTADO_LEDS: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		
		SAIDA_OPERACAO_DISPLAY: OUT STD_LOGIC_VECTOR (0 TO 6);	
		
		PUSH_RESULTADO: IN STD_LOGIC;
		PUSH_OPERACAO: IN STD_LOGIC;
		CLOCK: IN STD_LOGIC;
		LED_REFERENCIA: OUT STD_LOGIC
		
	);
END PROJETO;

ARCHITECTURE MODELO OF PROJETO IS 

CONSTANT CLOCK_FREE : INTEGER := 50e6;
SIGNAL TICKS : INTEGER := 0;
SIGNAL SEGUNDOS: INTEGER := 0;

SIGNAL OPERACAO: INTEGER := 1;

-- GUARDANDO RESULTADOS
SIGNAL RESULTADO_ARI: INTEGER := 0;
SIGNAL RESULTADO_LOG: STD_LOGIC_VECTOR (0 DOWNTO 5);

-- TRANSFORMANDO ENTRADA EM VALOR NÚMERICO
SIGNAL VALOR_1: INTEGER := TO_INTEGER(UNSIGNED(ENTRADA_1)); 
SIGNAL VALOR_2: INTEGER := TO_INTEGER(UNSIGNED(ENTRADA_2));


BEGIN
	
	PROCESS (CLOCK) IS
	BEGIN
	
		IF RISING_EDGE(CLOCK) THEN -- NA BORDA DO CLOCK
			IF TICKS = CLOCK_FREE - 1 THEN
				TICKS <= 0;
				-- CONTADOR DE TICKS
				IF SEGUNDOS = 3 THEN -- VAI aGIR APENAS QUANDO BATER 3S 
					SEGUNDOS <= 0;
					LED_REFERENCIA <= '1';
					CASE OPERACAO IS
						
						WHEN 1 => -- SOMA
						
							IF SINAL_1 = '0' THEN
								 VALOR_1 <= -VALOR_1;
							END IF;
							IF SINAL_2 = '0' THEN
								 VALOR_2 <= -VALOR_2;
							END IF;
							
							RESULTADO_ARI <= VALOR_1 + VALOR_2;
							
						WHEN 2 => -- ADIÇÃO
							
							IF SINAL_1 = '0' THEN
								 VALOR_1 <= -VALOR_1;
							END IF;
							IF SINAL_2 = '0' THEN
								 VALOR_2 <= -VALOR_2;
							END IF;
							
							RESULTADO_ARI <= VALOR_1 - VALOR_2;
						
						WHEN 3 => -- E
							
							RESULTADO_LOG <= ENTRADA_1 AND ENTRADA_2;
							
						WHEN 4 => -- OU
							
							RESULTADO_LOG <= ENTRADA_1 OR ENTRADA_2;
							
						WHEN 5 => -- OU EXCLUSUVIO
							
							RESULTADO_LOG <= ENTRADA_1 XOR ENTRADA_2;
							
						WHEN OTHERS => -- COMPLEMENTO	
							 
							RESULTADO_LOG <= NOT ENTRADA_1;
							
					END CASE;
					
				ELSE
					SEGUNDOS <= SEGUNDOS + 1;
					LED_REFERENCIA <= '0';
				END IF;
				
			ELSE
				TICKS <= ticks + 1;
			END IF;
		END IF;
		
		IF PUSH_OPERACAO = '0' THEN -- INCREMENTO DA OPERAÇÃO
			
			OPERACAO <= OPERACAO + 1;
			
			IF OPERACAO = 7 THEN
				OPERACAO <= 1;
			END IF;
			
			TICKS <= 0;
			SEGUNDOS <= 0;
			OPERACAO <= 1;
			RESULTADO_DISPLAY_1 <= "1111111";
			RESULTADO_DISPLAY_2 <= "1111111";
			RESULTADO_DISPLAY_3 <= "1111111";
			LED_REFERENCIA <= '1';
			RESULTADO_ARI <= 0;
			RESULTADO_LOG <= "1111111";
			
			-- A cada troca de operação ele reseta tudo
			
		END IF;
		
		IF PUSH_RESULTADO = '0' THEN -- MOSTRAR O RESULTADO
			IF OPERACAO < 3 THEN
					-- OPERAÇÕES ARITMETICAS
			ELSE
			      -- OPERAÇÕES LÓGICAS
			END IF;
		END IF;
		
		
	END PROCESS;

	SAIDA_OPERACAO_DISPLAY <=  "1000000" when OPERACAO = 0 else
										"1111001" when OPERACAO = 1 else
										"0100100" when OPERACAO = 2 else
										"0110000" when OPERACAO = 3 else	
										"0011001" when OPERACAO = 4 else
										"0010010" when OPERACAO = 5 else
										"0000010" when OPERACAO = 6 else
										"1111000" when OPERACAO = 7 else
										"0000000" when OPERACAO = 8 else
										"0010000" when OPERACAO = 9 else	
										"0100000" when OPERACAO = 10 else
										"0000011" when OPERACAO = 11 else
										"1000110" when OPERACAO = 12 else
										"0100001" when OPERACAO = 13 else
										"0000110" when OPERACAO = 14 else
										"0001110" when OPERACAO = 15;
		
	
END MODELO;