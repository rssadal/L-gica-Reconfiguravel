LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;


ENTITY PROJETO IS
	PORT(
		
		ENTRADA_1: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		ENTRADA_2: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		
		SAIDA_RESULTADO: OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
		SAIDA_OPERACAO_DISPLAY: OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
		
		SAIDA_OPERACAO_LEDS: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		
		PUSH_RESULTADO: IN STD_LOGIC;
		PUSH_OPERACAO: IN STD_LOGIC;
		RESET: IN STD_LOGIC;
		CLOCK: IN STD_LOGIC
	);
END PROJETO;

ARCHITECTURE MODELO OF PROJETO IS 

CONSTANT CLOCK_FREE : INTEGER := 50e6;
SIGNAL TICKS : INTEGER := 0;
SIGNAL SEGUNDOS: INTEGER := 0;
SIGNAL OPERACAO: INTEGER := 1;
SIGNAL RESULTADO: STD_LOGIC_VECTOR (3 DOWNTO 0);

BEGIN
	
	PROCESS (CLOCK) IS
	BEGIN
	
		IF RISING_EDGE(CLOCK) THEN -- NA BORDA DO CLOCK
			IF TICKS = CLOCK_FREE - 1 THEN
				TICKS <= 0;
				-- CONTADOR DE TICKS
				IF SEGUNDOS = 1 THEN -- VAI aGIR APENAS QUANDO BATER 1S 
					SEGUNDOS <= 0;
					
					CASE OPERACAO IS
						
						WHEN 1 => -- SOMA
							RESULTADO <= std_logic_vector(unsigned(ENTRADA_1) + unsigned(ENTRADA_2)));
						WHEN 2 => -- ADIÇÃO
							RESULTADO <= std_logic_vector(unsigned(ENTRADA_1) - unsigned(ENTRADA_2)));
						WHEN 3 => -- E
							RESULTADO <= ENTRADA_1 AND ENTRADA_2
						WHEN 4 => -- OU
							RESULTADO <= ENTRADA_1 OR ENTRADA_2
						WHEN 5 => -- OU EXCLUSUVIO
							RESULTADO <= ENTRADA_1 XOR ENTRADA_2
						WHEN 6 => -- COMPLEMENTO	
							RESULTADO <= ENTRADA_1 NOT ENTRADA_2 
					END CASE;
					
				ELSE
					SEGUNDOS <= SEGUNDOS + 1;
				END IF;
				
			ELSE
				TICKS <= ticks + 1;
			END IF;
		END IF;
		
		IF RESET = '0' THEN
			TICKS <= 0;
			SEGUNDOS <= 0;
			OPERACAO <= 1;
			-- RESETAR TUDO 
		END IF;
		
		IF PUSH_OPERACAO = '0' THEN -- INCREMENTO DA OPERAÇÃO
			OPERACAO <= OPERACAO + 1;
			IF OPERACAO = 6
				OPERACAO <= 1;
			END IF;
		END IF;

	END PROCESS;

END MODELO;